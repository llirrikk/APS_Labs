module rom256_32 (         // создать блок с именем rom256_32
  input   [31:0]   A,      // 32-битный адресный вход
  output  [255:0]  RD      // 256-битный выход считанных данных
);

  reg [31:0] ROM [0:255];   // создать память с 256-ю 32-битными ячейками


  initial $readmemb("mem.txt", RAM);  // поместить при запуске микросхемы в
                                      // память RAM содержимое файла mem.txt

   

  assign RD = ROM[A];   // реализация первого порта на чтение

endmodule                 //  конец описания модуля

