module rom32_8 (          // создать блок с именем rom32_8
  input   [7:0]   A,      // 8-битный адресный вход
  output  [31:0]  RD      // 32-битный выход считанных данных
);

  reg [7:0] ROM [0:31];   // создать память с 32-ю 8-битными ячейками


  initial $readmemb("mem.txt", ROM);  // поместить при запуске микросхемы в
                                      // память ROM содержимое файла mem.txt

   

  assign RD = ROM[A];   // реализация первого порта на чтение

endmodule                 //  конец описания модуля

